library IEEE;
use IEEE.STD_LOGIC_1164.all;

package MyTypes is

    type states is (idle, start_bit, stop_bit, data_bits, reset_check);

end MyTypes;

package body MyTypes is
end MyTypes;